CIRCUIT D:\Documents and Settings\sicard\Mes documents\software\Microwind\microwind35\examples\inverter\cmos.MSK
*
* IC Technology: CMOS 45nm - HighK/Metal/Strain - 8 Metal copper
*
VDD 1 0 DC 1.00
VA 5 0 DC 0 PULSE(0.00 1.00 0.95N 0.05N 0.05N 0.95N 2.00N)
*
* List of nodes
* "nA" corresponds to n�3
* "A" corresponds to n�5
*
* MOS devices
MN1 0 5 3 0 N1  W= 0.20U L= 0.04U
MP1 3 5 1 1 P1  W= 0.20U L= 0.04U
*
C2 1 0  0.148fF
C3 3 0  0.180fF
C5 5 0  0.072fF
*
* n-MOS Model 3 :
* low leakage
.MODEL N1 NMOS LEVEL=3 VTO=0.18 UO=160.000 TOX= 3.5E-9
+LD =0.005U THETA=0.300 GAMMA=0.400
+PHI=0.150 KAPPA=0.350 VMAX=180.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* p-MOS Model 3:
* low leakage
.MODEL P1 PMOS LEVEL=3 VTO=-0.15 UO=120.000 TOX= 3.5E-9
+LD =0.005U THETA=0.300 GAMMA=0.400
+PHI=0.150 KAPPA=0.350 VMAX=180.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
* (Winspice)
.options temp=27.0
.control
tran 0.1N 1.00N
print  V(3) V(5) > out.txt
plot  V(3) V(5)
.endc
.END
