CIRCUIT D:\Documents and Settings\sicard\Mes documents\software\Microwind\microwind35\examples\adders\halfAdder.MSK
*
* IC Technology: CMOS 45nm - HighK/Metal - 3rd generation Strain - 8 Metal copper
*
VDD 1 0 DC 1.00
VA 9 0 DC 0 PULSE(0.00 1.00 1.98N 0.02N 0.02N 1.98N 4.00N)
VB 11 0 DC 0 PULSE(0.00 1.00 0.98N 0.02N 0.02N 0.98N 2.00N)
*
* List of nodes
* " xor2_Sum" corresponds to n�3
* "N4" corresponds to n�4
* "N5" corresponds to n�5
* " and2_Carry" corresponds to n�7
* "N8" corresponds to n�8
* "A" corresponds to n�9
* "B" corresponds to n�11
*
* MOS devices
MN1 0 4 3 0 N1  W= 0.22U L= 0.04U
MN2 9 11 4 0 N1  W= 0.14U L= 0.04U
MN3 0 9 5 0 N1  W= 0.08U L= 0.04U
MN4 0 8 7 0 N1  W= 0.08U L= 0.04U
MN5 10 9 8 0 N1  W= 0.08U L= 0.04U
MN6 0 11 10 0 N1  W= 0.08U L= 0.04U
MP1 1 4 3 1 P1  W= 0.24U L= 0.04U
MP2 5 11 4 1 P1  W= 0.24U L= 0.04U
MP3 1 9 5 1 P1  W= 0.24U L= 0.04U
MP4 1 8 7 1 P1  W= 0.24U L= 0.04U
MP5 8 9 1 1 P1  W= 0.24U L= 0.04U
MP6 1 11 8 1 P1  W= 0.24U L= 0.04U
*
C2 1 0  1.092fF
C3 3 0  0.535fF
C4 4 0  0.286fF
C5 5 0  0.163fF
C7 7 0  0.410fF
C8 8 0  0.289fF
C9 9 0  0.535fF
C10 10 0  0.019fF
C11 11 0  0.452fF
*
*
* n-MOS BSIM4 :
* low leakage
.MODEL N1 NMOS LEVEL=14 VTHO=0.24 U0=0.034 TOXE= 2.0E-9 LINT=0.000U 
+K1 =0.750 K2=0.100 DVT0=2.300
+DVT1=0.540 LPE0=2.200e-9 ETA0=0.080
+NFACTOR=  0.5 UA=6.300e-15
+WINT=0.020U UC=-0.047e-15 PSCBE1=230.000e6
+KT1=-0.060 UTE=-1.800
+XJ=0.150U NDEP=170.000e15 PCLM=1.100
+VSAT=100000.000 VOFF=0.000
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* p-MOS BSIM4:
* low leakage
.MODEL P1 PMOS LEVEL=14 VTHO=-0.15 U0=0.024 TOXE= 2.0E-9 LINT=0.000U 
+K1 =0.500 K2=0.100 DVT0=2.300
+DVT1=0.540 LPE0=2.200e-9 ETA0=0.080
+NFACTOR=  0.4 UA=9.500e-15
+WINT=0.020U UC=-0.047e-15 PSCBE1=230.000e6
+KT1=-0.060 UTE=-1.800
+XJ=0.150U NDEP=170.000e15 PCLM=0.700
+VSAT=60000.000 VOFF=0.000
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* Transient analysis
*
* (Winspice)
.options temp=27.0
.control
tran 0.1N 5.00N
print  V(11) V(9) V(7) V(3) > out.txt
plot  V(11) V(9) V(7) V(3)
.endc
.END
