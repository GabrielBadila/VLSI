// DSCH 3.5
// 31/08/2009 09:08:27
// D:\Documents and Settings\sicard\Mes documents\software\Dsch\Dsch35\dsch35 full\examples\test\input_order.sch

module input_order( C,Bs,A);
 input C,Bs,A;
 wire ;
endmodule

// Simulation parameters in Verilog Format
always
#200 C=~C;
#400 B>=~B>;
#800 A=~A;

// Simulation parameters
// C CLK 1 1
// B> CLK 2 2
// A CLK 4 4
